-- ====================================================================
--
--	File Name:		Idecode.vhd
--	Description:	Idecode module (implements the register file for the MIPS computer)
--
--
--	Date:			30/05/2018
--	Designers:		Maor Assayag, Refael Shetrit
--
-- ====================================================================

-- libraries decleration
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

 -- entity Definition
ENTITY Idecode IS
	  PORT(	read_data_1	: OUT 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
			read_data_2	: OUT 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
			old_Instruction : IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
			Instruction : IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
			read_data 	: IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
			ALU_result	: IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
			RegWrite 	: IN 	STD_LOGIC;
			MemtoReg 	: IN 	STD_LOGIC;
			RegDst 		: IN 	STD_LOGIC;
			Sign_extend : OUT 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
			clock,reset,button_GPIO	: IN 	STD_LOGIC ;
			LO_1    			    :     out  std_logic_vector (6 downto 0);
			LO_2    				 :     out  std_logic_vector (6 downto 0);
			HI_1    				 :     out  std_logic_vector (6 downto 0);
			HI_2   				 :     out  std_logic_vector (6 downto 0));
END Idecode;

 -- Architecture Definition
ARCHITECTURE behavior OF Idecode IS
COMPONENT display_7_segment
    port (
    	q        : in std_logic_vector (7 downto 0);
    	segment1 : out std_logic_vector (6 downto 0);
      segment2 : out std_logic_vector (6 downto 0));
end COMPONENT;

COMPONENT Counter  port (
	clk,enable : in std_logic;
	q          : out std_logic_vector (7 downto 0));
end COMPONENT;
TYPE register_file IS ARRAY ( 0 TO 31 ) OF STD_LOGIC_VECTOR( 31 DOWNTO 0 );

	SIGNAL register_array				: register_file;
	SIGNAL write_register_address 		: STD_LOGIC_VECTOR( 4 DOWNTO 0 );
	SIGNAL write_data					      : STD_LOGIC_VECTOR( 31 DOWNTO 0 );
	SIGNAL read_register_1_address		: STD_LOGIC_VECTOR( 4 DOWNTO 0 );
	SIGNAL read_register_2_address		: STD_LOGIC_VECTOR( 4 DOWNTO 0 );
	SIGNAL write_register_address_1		: STD_LOGIC_VECTOR( 4 DOWNTO 0 );
	SIGNAL write_register_address_0		: STD_LOGIC_VECTOR( 4 DOWNTO 0 );
	SIGNAL Instruction_immediate_value	: STD_LOGIC_VECTOR( 15 DOWNTO 0 );
	SIGNAL en_7_seg          :     STD_LOGIC:= '0';
	SIGNAL i          :     integer := 0;
   SIGNAL q                 :     STD_LOGIC_VECTOR ( 7 DOWNTO 0 );
   SIGNAL memread                 :     STD_LOGIC_VECTOR ( 31 DOWNTO 0 );



BEGIN
----------------------------------------
		read_register_1_address 	<= Instruction( 25 DOWNTO 21 );
   	read_register_2_address 	<= Instruction( 20 DOWNTO 16 );
   	write_register_address_1	<= old_Instruction( 15 DOWNTO 11 );
   	write_register_address_0 	<= old_Instruction( 20 DOWNTO 16 );
   	Instruction_immediate_value <= Instruction( 15 DOWNTO 0 );
					-- Read Register 1 Operation
	read_data_1 <= write_data
	WHEN (write_register_address = read_register_1_address) and RegWrite = '1'
	ELSE register_array(
			      CONV_INTEGER( read_register_1_address ) );
					-- Read Register 2 Operation
	read_data_2 <= write_data
	WHEN write_register_address = read_register_2_address  and RegWrite = '1'
	ELSE register_array(
			      CONV_INTEGER( read_register_2_address ) );
					-- Mux for Register Write Address
    	write_register_address <= write_register_address_1
			WHEN RegDst = '1'  			ELSE write_register_address_0;
					-- Mux to bypass data memory for Rformat instructions
	write_data <= ALU_result( 31 DOWNTO 0 )
			WHEN ( MemtoReg = '0' ) 	ELSE read_data;
					-- Sign Extend 16-bits to 32-bits
    	Sign_extend <= X"0000" & Instruction_immediate_value
		WHEN Instruction_immediate_value(15) = '0'
		ELSE	X"FFFF" & Instruction_immediate_value;

PROCESS (clock, write_register_address, RegWrite, write_data)
	variable zero : STD_LOGIC_VECTOR (31 downto 0) := (others => '0');
	BEGIN
		IF rising_edge(clock) THEN
		IF reset = '1' THEN
					-- Initial register values on reset are register = reg#
					-- use loop to automatically generate reset logic
					-- for all registers
			FOR i IN 0 TO 31 LOOP
				register_array(i) <= zero;
 			END LOOP;
					-- Write back to register - don't write to register 0
  		ELSIF RegWrite = '1' AND write_register_address /= 0 THEN
		      register_array( CONV_INTEGER( write_register_address)) <= write_data;
		END IF;
		END IF;
	END PROCESS;
----------------------------------------







counter_en:process (button_GPIO)
						begin
								if (rising_edge(button_GPIO)) then
										en_7_seg <= '1';
							 end if;
						end process;


-------------------------------        display
Counter_unit : Counter
			PORT MAP (
					clk => clock,
					enable => en_7_seg,
					q => q
			);



display7 : process
begin
wait until q(1)'event and q(1) = '1';
		if i < 8 then
			i <= i+1;
		end if;
end process;

memread <=   register_array(i+ 14) when i < 8 else (31 downto 0 =>'0') ;
convert_7_segment_1: display_7_segment port map (memread( 7 downto 0),LO_1, LO_2);
convert_7_segment_2: display_7_segment port map (memread(15 downto 8),HI_1,HI_2);






END behavior;

--EndOfFile
